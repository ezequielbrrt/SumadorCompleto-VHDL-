module sumadorcompleto ( 
	x,
	y,
	z,
	a,
	s
	) ;

input  x;
input  y;
input  z;
inout  a;
inout  s;
